library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity instr_decoder is 
end entity;

architecture behav of instr_decoder is
      
begin
    
    
    
end architecture behav;

