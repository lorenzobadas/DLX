library ieee;
use ieee.std_logic_1164.all;
package instructions_pkg is
-- MANDATORY INSTRUCTIONS
    -- OPCODE FIELD
    constant opcode_j:       std_logic_vector(5 downto 0) := "000010";       -- 0x02
    constant opcode_jal:     std_logic_vector(5 downto 0) := "000011";       -- 0x03
    constant opcode_beqz:    std_logic_vector(5 downto 0) := "000100";       -- 0x04
    constant opcode_bnez:    std_logic_vector(5 downto 0) := "000101";       -- 0x05
    constant opcode_addi:    std_logic_vector(5 downto 0) := "001000";       -- 0x08
    constant opcode_subi:    std_logic_vector(5 downto 0) := "001010";       -- 0x0a
    constant opcode_andi:    std_logic_vector(5 downto 0) := "001100";       -- 0x0c
    constant opcode_ori:     std_logic_vector(5 downto 0) := "001101";       -- 0x0d
    constant opcode_xori:    std_logic_vector(5 downto 0) := "001110";       -- 0x0e
    constant opcode_slli:    std_logic_vector(5 downto 0) := "010100";       -- 0x14
    constant opcode_nop:     std_logic_vector(5 downto 0) := "010101";       -- 0x15
    constant opcode_srli:    std_logic_vector(5 downto 0) := "010110";       -- 0x16
    constant opcode_snei:    std_logic_vector(5 downto 0) := "011001";       -- 0x19
    constant opcode_slei:    std_logic_vector(5 downto 0) := "011100";       -- 0x1c
    constant opcode_sgei:    std_logic_vector(5 downto 0) := "011101";       -- 0x1d
    constant opcode_lw:      std_logic_vector(5 downto 0) := "100011";       -- 0x23
    constant opcode_sw:      std_logic_vector(5 downto 0) := "101011";       -- 0x2b
    constant opcode_sll:     std_logic_vector(5 downto 0) := "000000";       -- 0x0
    constant opcode_srl:     std_logic_vector(5 downto 0) := "000000";       -- 0x0
    constant opcode_add:     std_logic_vector(5 downto 0) := "000000";       -- 0x0
    constant opcode_sub:     std_logic_vector(5 downto 0) := "000000";       -- 0x0
    constant opcode_and:     std_logic_vector(5 downto 0) := "000000";       -- 0x0
    constant opcode_or:      std_logic_vector(5 downto 0) := "000000";       -- 0x0
    constant opcode_xor:     std_logic_vector(5 downto 0) := "000000";       -- 0x0
    constant opcode_sne:     std_logic_vector(5 downto 0) := "000000";       -- 0x0
    constant opcode_sle:     std_logic_vector(5 downto 0) := "000000";       -- 0x0
    constant opcode_sge:     std_logic_vector(5 downto 0) := "000000";       -- 0x0

    -- FUNC FIELD
    constant func_sll:       std_logic_vector(10 downto 0) := "00000000100"; -- 0x04
    constant func_srl:       std_logic_vector(10 downto 0) := "00000000110"; -- 0x06
    constant func_add:       std_logic_vector(10 downto 0) := "00000100000"; -- 0x20
    constant func_sub:       std_logic_vector(10 downto 0) := "00000100010"; -- 0x22
    constant func_and:       std_logic_vector(10 downto 0) := "00000100100"; -- 0x24
    constant func_or:        std_logic_vector(10 downto 0) := "00000100101"; -- 0x25
    constant func_xor:       std_logic_vector(10 downto 0) := "00000100110"; -- 0x26
    constant func_sne:       std_logic_vector(10 downto 0) := "00000101001"; -- 0x29
    constant func_sle:       std_logic_vector(10 downto 0) := "00000101100"; -- 0x2c
    constant func_sge:       std_logic_vector(10 downto 0) := "00000101101"; -- 0x2d

-- OPTIONAL INSTRUCTIONS
    -- OPCODE FIELD
    constant opcode_bfpt:    std_logic_vector(5 downto 0) := "000110";       -- 0x06
    constant opcode_bfpf:    std_logic_vector(5 downto 0) := "000111";       -- 0x07
    constant opcode_addui:   std_logic_vector(5 downto 0) := "001001";       -- 0x09
    constant opcode_subui:   std_logic_vector(5 downto 0) := "001011";       -- 0x0b
    constant opcode_lhi:     std_logic_vector(5 downto 0) := "001111";       -- 0x0f
    constant opcode_rfe:     std_logic_vector(5 downto 0) := "010000";       -- 0x10
    constant opcode_trap:    std_logic_vector(5 downto 0) := "010001";       -- 0x11
    constant opcode_jr:      std_logic_vector(5 downto 0) := "010010";       -- 0x12
    constant opcode_jalr:    std_logic_vector(5 downto 0) := "010011";       -- 0x13
    constant opcode_srai:    std_logic_vector(5 downto 0) := "010111";       -- 0x17
    constant opcode_seqi:    std_logic_vector(5 downto 0) := "011000";       -- 0x18
    constant opcode_slti:    std_logic_vector(5 downto 0) := "011010";       -- 0x1a
    constant opcode_sgti:    std_logic_vector(5 downto 0) := "011011";       -- 0x1b
    constant opcode_lb:      std_logic_vector(5 downto 0) := "100000";       -- 0x20
    constant opcode_lh:      std_logic_vector(5 downto 0) := "100001";       -- 0x21
    constant opcode_lbu:     std_logic_vector(5 downto 0) := "100100";       -- 0x24
    constant opcode_lhu:     std_logic_vector(5 downto 0) := "100101";       -- 0x25
    constant opcode_lf:      std_logic_vector(5 downto 0) := "100110";       -- 0x26
    constant opcode_ld:      std_logic_vector(5 downto 0) := "100111";       -- 0x27
    constant opcode_sb:      std_logic_vector(5 downto 0) := "101000";       -- 0x28
    constant opcode_sh:      std_logic_vector(5 downto 0) := "101001";       -- 0x29
    constant opcode_sf:      std_logic_vector(5 downto 0) := "101110";       -- 0x2e
    constant opcode_sd:      std_logic_vector(5 downto 0) := "101111";       -- 0x2f
    constant opcode_itlb:    std_logic_vector(5 downto 0) := "111000";       -- 0x38
    constant opcode_sltui:   std_logic_vector(5 downto 0) := "111010";       -- 0x3a
    constant opcode_sgtui:   std_logic_vector(5 downto 0) := "111011";       -- 0x3b
    constant opcode_sleui:   std_logic_vector(5 downto 0) := "111100";       -- 0x3c
    constant opcode_sgeui:   std_logic_vector(5 downto 0) := "111101";       -- 0x3d
    constant opcode_sra:     std_logic_vector(5 downto 0) := "000000";       -- 0x0
    constant opcode_addu:    std_logic_vector(5 downto 0) := "000000";       -- 0x0
    constant opcode_subu:    std_logic_vector(5 downto 0) := "000000";       -- 0x0
    constant opcode_seq:     std_logic_vector(5 downto 0) := "000000";       -- 0x0
    constant opcode_slt:     std_logic_vector(5 downto 0) := "000000";       -- 0x0
    constant opcode_sgt:     std_logic_vector(5 downto 0) := "000000";       -- 0x0
    constant opcode_movi2s:  std_logic_vector(5 downto 0) := "000000";       -- 0x0
    constant opcode_movs2i:  std_logic_vector(5 downto 0) := "000000";       -- 0x0
    constant opcode_movf:    std_logic_vector(5 downto 0) := "000000";       -- 0x0
    constant opcode_movd:    std_logic_vector(5 downto 0) := "000000";       -- 0x0
    constant opcode_movfp2i: std_logic_vector(5 downto 0) := "000000";       -- 0x0
    constant opcode_movi2fp: std_logic_vector(5 downto 0) := "000000";       -- 0x0
    constant opcode_movi2t:  std_logic_vector(5 downto 0) := "000000";       -- 0x0
    constant opcode_movt2i:  std_logic_vector(5 downto 0) := "000000";       -- 0x0
    constant opcode_sltu:    std_logic_vector(5 downto 0) := "000000";       -- 0x0
    constant opcode_sgtu:    std_logic_vector(5 downto 0) := "000000";       -- 0x0
    constant opcode_sleu:    std_logic_vector(5 downto 0) := "000000";       -- 0x0
    constant opcode_sgeu:    std_logic_vector(5 downto 0) := "000000";       -- 0x0
    constant opcode_addf:    std_logic_vector(5 downto 0) := "000100";       -- 0x4
    constant opcode_subf:    std_logic_vector(5 downto 0) := "000100";       -- 0x4
    constant opcode_multf:   std_logic_vector(5 downto 0) := "000100";       -- 0x4
    constant opcode_divf:    std_logic_vector(5 downto 0) := "000100";       -- 0x4
    constant opcode_addd:    std_logic_vector(5 downto 0) := "000100";       -- 0x4
    constant opcode_subd:    std_logic_vector(5 downto 0) := "000100";       -- 0x4
    constant opcode_multd:   std_logic_vector(5 downto 0) := "000100";       -- 0x4
    constant opcode_divd:    std_logic_vector(5 downto 0) := "000100";       -- 0x4
    constant opcode_cvtf2d:  std_logic_vector(5 downto 0) := "000100";       -- 0x4
    constant opcode_cvtf2i:  std_logic_vector(5 downto 0) := "000100";       -- 0x4
    constant opcode_cvtd2f:  std_logic_vector(5 downto 0) := "000100";       -- 0x4
    constant opcode_cvtd2i:  std_logic_vector(5 downto 0) := "000100";       -- 0x4
    constant opcode_cvti2f:  std_logic_vector(5 downto 0) := "000100";       -- 0x4
    constant opcode_cvti2d:  std_logic_vector(5 downto 0) := "000100";       -- 0x4
    constant opcode_mult:    std_logic_vector(5 downto 0) := "000100";       -- 0x4
    constant opcode_div:     std_logic_vector(5 downto 0) := "000100";       -- 0x4
    constant opcode_eqf:     std_logic_vector(5 downto 0) := "000100";       -- 0x4
    constant opcode_nef:     std_logic_vector(5 downto 0) := "000100";       -- 0x4
    constant opcode_ltf:     std_logic_vector(5 downto 0) := "000100";       -- 0x4
    constant opcode_gtf:     std_logic_vector(5 downto 0) := "000100";       -- 0x4
    constant opcode_lef:     std_logic_vector(5 downto 0) := "000100";       -- 0x4
    constant opcode_gef:     std_logic_vector(5 downto 0) := "000100";       -- 0x4
    constant opcode_multu:   std_logic_vector(5 downto 0) := "000100";       -- 0x4
    constant opcode_divu:    std_logic_vector(5 downto 0) := "000100";       -- 0x4
    constant opcode_eqd:     std_logic_vector(5 downto 0) := "000100";       -- 0x4
    constant opcode_ned:     std_logic_vector(5 downto 0) := "000100";       -- 0x4
    constant opcode_ltd:     std_logic_vector(5 downto 0) := "000100";       -- 0x4
    constant opcode_gtd:     std_logic_vector(5 downto 0) := "000100";       -- 0x4
    constant opcode_led:     std_logic_vector(5 downto 0) := "000100";       -- 0x4
    constant opcode_ged:     std_logic_vector(5 downto 0) := "000100";       -- 0x4

    -- FUNC FIELD
    constant func_sra:       std_logic_vector(10 downto 0) := "00000000111"; -- 0x07
    constant func_addu:      std_logic_vector(10 downto 0) := "00000100001"; -- 0x21
    constant func_subu:      std_logic_vector(10 downto 0) := "00000100011"; -- 0x23
    constant func_seq:       std_logic_vector(10 downto 0) := "00000101000"; -- 0x28
    constant func_slt:       std_logic_vector(10 downto 0) := "00000101010"; -- 0x2a
    constant func_sgt:       std_logic_vector(10 downto 0) := "00000101011"; -- 0x2b
    constant func_movi2s:    std_logic_vector(10 downto 0) := "00000110000"; -- 0x30
    constant func_movs2i:    std_logic_vector(10 downto 0) := "00000110001"; -- 0x31
    constant func_movf:      std_logic_vector(10 downto 0) := "00000110010"; -- 0x32
    constant func_movd:      std_logic_vector(10 downto 0) := "00000110011"; -- 0x33
    constant func_movfp2i:   std_logic_vector(10 downto 0) := "00000110100"; -- 0x34
    constant func_movi2fp:   std_logic_vector(10 downto 0) := "00000110101"; -- 0x35
    constant func_movi2t:    std_logic_vector(10 downto 0) := "00000110110"; -- 0x36
    constant func_movt2i:    std_logic_vector(10 downto 0) := "00000110111"; -- 0x37
    constant func_sltu:      std_logic_vector(10 downto 0) := "00000111010"; -- 0x3a
    constant func_sgtu:      std_logic_vector(10 downto 0) := "00000111011"; -- 0x3b
    constant func_sleu:      std_logic_vector(10 downto 0) := "00000111100"; -- 0x3c
    constant func_sgeu:      std_logic_vector(10 downto 0) := "00000111101"; -- 0x3d
    constant func_addf:      std_logic_vector(10 downto 0) := "00000000000"; -- 0x00
    constant func_subf:      std_logic_vector(10 downto 0) := "00000000001"; -- 0x01
    constant func_multf:     std_logic_vector(10 downto 0) := "00000000010"; -- 0x02
    constant func_divf:      std_logic_vector(10 downto 0) := "00000000011"; -- 0x03
    constant func_addd:      std_logic_vector(10 downto 0) := "00000000100"; -- 0x04
    constant func_subd:      std_logic_vector(10 downto 0) := "00000000101"; -- 0x05
    constant func_multd:     std_logic_vector(10 downto 0) := "00000000110"; -- 0x06
    constant func_divd:      std_logic_vector(10 downto 0) := "00000000111"; -- 0x07
    constant func_cvtf2d:    std_logic_vector(10 downto 0) := "00000001000"; -- 0x08
    constant func_cvtf2i:    std_logic_vector(10 downto 0) := "00000001001"; -- 0x09
    constant func_cvtd2f:    std_logic_vector(10 downto 0) := "00000001010"; -- 0x0a
    constant func_cvtd2i:    std_logic_vector(10 downto 0) := "00000001011"; -- 0x0b
    constant func_cvti2f:    std_logic_vector(10 downto 0) := "00000001100"; -- 0x0c
    constant func_cvti2d:    std_logic_vector(10 downto 0) := "00000001101"; -- 0x0d
    constant func_mult:      std_logic_vector(10 downto 0) := "00000001110"; -- 0x0e
    constant func_div:       std_logic_vector(10 downto 0) := "00000001111"; -- 0x0f
    constant func_eqf:       std_logic_vector(10 downto 0) := "00000010000"; -- 0x10
    constant func_nef:       std_logic_vector(10 downto 0) := "00000010001"; -- 0x11
    constant func_ltf:       std_logic_vector(10 downto 0) := "00000010010"; -- 0x12
    constant func_gtf:       std_logic_vector(10 downto 0) := "00000010011"; -- 0x13
    constant func_lef:       std_logic_vector(10 downto 0) := "00000010100"; -- 0x14
    constant func_gef:       std_logic_vector(10 downto 0) := "00000010101"; -- 0x15
    constant func_multu:     std_logic_vector(10 downto 0) := "00000010110"; -- 0x16
    constant func_divu:      std_logic_vector(10 downto 0) := "00000010111"; -- 0x17
    constant func_eqd:       std_logic_vector(10 downto 0) := "00000011000"; -- 0x18
    constant func_ned:       std_logic_vector(10 downto 0) := "00000011001"; -- 0x19
    constant func_ltd:       std_logic_vector(10 downto 0) := "00000011010"; -- 0x1a
    constant func_gtd:       std_logic_vector(10 downto 0) := "00000011011"; -- 0x1b
    constant func_led:       std_logic_vector(10 downto 0) := "00000011100"; -- 0x1c
    constant func_ged:       std_logic_vector(10 downto 0) := "00000011101"; -- 0x1d

end instructions_pkg;
