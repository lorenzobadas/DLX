library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity mem_wb_regs is
    generic(
        nbit : integer := 32
    );
    port (
        clk_i       : in  std_logic;
        reset_i     : in  std_logic;
        aluout_i    : in  std_logic_vector(nbit-1 downto 0);
        dout_i       : in  std_logic_vector(nbit-1 downto 0);
        rdest_i     : in  std_logic_vector(4 downto 0);
        aluout_o    : out std_logic_vector(nbit-1 downto 0);
        dout_o       : out std_logic_vector(nbit-1 downto 0);
        rdest_o     : out std_logic_vector(4 downto 0);
        -- Control signals
        memToReg_i  : in std_logic;
        regWrite_i  : in std_logic;
        memToReg_o  : out std_logic;
        regWrite_o  : out std_logic
    );
end mem_wb_regs;

architecture behav of mem_wb_regs is
begin
    process(clk_i, reset_i)
    begin
        if reset_i = '1' then
            aluout_o <= (others => '0');
            dout_o <= (others => '0');
            rdest_o <= (others => '0');
            memToReg_o <= '0';
            regWrite_o <= '0';
        elsif rising_edge(clk_i) then
            aluout_o <= aluout_i;
            dout_o <= dout_i;
            rdest_o <= rdest_i;
            memToReg_o <= memToReg_i;
            regWrite_o <= regWrite_i;
        end if;
    end process;
end behav;
