��l i b r a r y   i e e e ;  
 u s e   i e e e . s t d _ l o g i c _ 1 1 6 4 . a l l ;  
 p a c k a g e   i n s t r u c t i o n s _ p k g   i s  
         - -   O P C O D E   F I E L D  
         c o n s t a n t   o p c o d e _ j :               s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 0 1 0 " ;               - -   0 x 0 2  
         c o n s t a n t   o p c o d e _ j a l :           s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 0 1 1 " ;               - -   0 x 0 3  
         c o n s t a n t   o p c o d e _ b e q z :         s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 1 0 0 " ;               - -   0 x 0 4  
         c o n s t a n t   o p c o d e _ b n e z :         s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 1 0 1 " ;               - -   0 x 0 5  
         c o n s t a n t   o p c o d e _ b f p t :         s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 1 1 0 " ;               - -   0 x 0 6  
         c o n s t a n t   o p c o d e _ b f p f :         s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 1 1 1 " ;               - -   0 x 0 7  
         c o n s t a n t   o p c o d e _ a d d i :         s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 1 0 0 0 " ;               - -   0 x 0 8  
         c o n s t a n t   o p c o d e _ a d d u i :       s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 1 0 0 1 " ;               - -   0 x 0 9  
         c o n s t a n t   o p c o d e _ s u b i :         s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 1 0 1 0 " ;               - -   0 x 0 a  
         c o n s t a n t   o p c o d e _ s u b u i :       s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 1 0 1 1 " ;               - -   0 x 0 b  
         c o n s t a n t   o p c o d e _ a n d i :         s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 1 1 0 0 " ;               - -   0 x 0 c  
         c o n s t a n t   o p c o d e _ o r i :           s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 1 1 0 1 " ;               - -   0 x 0 d  
         c o n s t a n t   o p c o d e _ x o r i :         s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 1 1 1 0 " ;               - -   0 x 0 e  
         c o n s t a n t   o p c o d e _ l h i :           s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 1 1 1 1 " ;               - -   0 x 0 f  
         c o n s t a n t   o p c o d e _ r f e :           s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 1 0 0 0 0 " ;               - -   0 x 1 0  
         c o n s t a n t   o p c o d e _ t r a p :         s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 1 0 0 0 1 " ;               - -   0 x 1 1  
         c o n s t a n t   o p c o d e _ j r :             s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 1 0 0 1 0 " ;               - -   0 x 1 2  
         c o n s t a n t   o p c o d e _ j a l r :         s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 1 0 0 1 1 " ;               - -   0 x 1 3  
         c o n s t a n t   o p c o d e _ s l l i :         s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 1 0 1 0 0 " ;               - -   0 x 1 4  
         c o n s t a n t   o p c o d e _ n o p :           s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 1 0 1 0 1 " ;               - -   0 x 1 5  
         c o n s t a n t   o p c o d e _ s r l i :         s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 1 0 1 1 0 " ;               - -   0 x 1 6  
         c o n s t a n t   o p c o d e _ s r a i :         s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 1 0 1 1 1 " ;               - -   0 x 1 7  
         c o n s t a n t   o p c o d e _ s e q i :         s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 1 1 0 0 0 " ;               - -   0 x 1 8  
         c o n s t a n t   o p c o d e _ s n e i :         s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 1 1 0 0 1 " ;               - -   0 x 1 9  
         c o n s t a n t   o p c o d e _ s l t i :         s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 1 1 0 1 0 " ;               - -   0 x 1 a  
         c o n s t a n t   o p c o d e _ s g t i :         s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 1 1 0 1 1 " ;               - -   0 x 1 b  
         c o n s t a n t   o p c o d e _ s l e i :         s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 1 1 1 0 0 " ;               - -   0 x 1 c  
         c o n s t a n t   o p c o d e _ s g e i :         s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 1 1 1 0 1 " ;               - -   0 x 1 d  
         c o n s t a n t   o p c o d e _ l b :             s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 1 0 0 0 0 0 " ;               - -   0 x 2 0  
         c o n s t a n t   o p c o d e _ l h :             s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 1 0 0 0 0 1 " ;               - -   0 x 2 1  
         c o n s t a n t   o p c o d e _ l w :             s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 1 0 0 0 1 1 " ;               - -   0 x 2 3  
         c o n s t a n t   o p c o d e _ l b u :           s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 1 0 0 1 0 0 " ;               - -   0 x 2 4  
         c o n s t a n t   o p c o d e _ l h u :           s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 1 0 0 1 0 1 " ;               - -   0 x 2 5  
         c o n s t a n t   o p c o d e _ l f :             s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 1 0 0 1 1 0 " ;               - -   0 x 2 6  
         c o n s t a n t   o p c o d e _ l d :             s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 1 0 0 1 1 1 " ;               - -   0 x 2 7  
         c o n s t a n t   o p c o d e _ s b :             s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 1 0 1 0 0 0 " ;               - -   0 x 2 8  
         c o n s t a n t   o p c o d e _ s h :             s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 1 0 1 0 0 1 " ;               - -   0 x 2 9  
         c o n s t a n t   o p c o d e _ s w :             s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 1 0 1 0 1 1 " ;               - -   0 x 2 b  
         c o n s t a n t   o p c o d e _ s f :             s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 1 0 1 1 1 0 " ;               - -   0 x 2 e  
         c o n s t a n t   o p c o d e _ s d :             s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 1 0 1 1 1 1 " ;               - -   0 x 2 f  
         c o n s t a n t   o p c o d e _ i t l b :         s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 1 1 1 0 0 0 " ;               - -   0 x 3 8  
         c o n s t a n t   o p c o d e _ s l t u i :       s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 1 1 1 0 1 0 " ;               - -   0 x 3 a  
         c o n s t a n t   o p c o d e _ s g t u i :       s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 1 1 1 0 1 1 " ;               - -   0 x 3 b  
         c o n s t a n t   o p c o d e _ s l e u i :       s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 1 1 1 1 0 0 " ;               - -   0 x 3 c  
         c o n s t a n t   o p c o d e _ s g e u i :       s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 1 1 1 1 0 1 " ;               - -   0 x 3 d  
         c o n s t a n t   o p c o d e _ s l l :           s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 0 0 0 " ;               - -   0 x 0  
         c o n s t a n t   o p c o d e _ s r l :           s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 0 0 0 " ;               - -   0 x 0  
         c o n s t a n t   o p c o d e _ s r a :           s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 0 0 0 " ;               - -   0 x 0  
         c o n s t a n t   o p c o d e _ a d d :           s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 0 0 0 " ;               - -   0 x 0  
         c o n s t a n t   o p c o d e _ a d d u :         s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 0 0 0 " ;               - -   0 x 0  
         c o n s t a n t   o p c o d e _ s u b :           s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 0 0 0 " ;               - -   0 x 0  
         c o n s t a n t   o p c o d e _ s u b u :         s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 0 0 0 " ;               - -   0 x 0  
         c o n s t a n t   o p c o d e _ a n d :           s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 0 0 0 " ;               - -   0 x 0  
         c o n s t a n t   o p c o d e _ o r :             s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 0 0 0 " ;               - -   0 x 0  
         c o n s t a n t   o p c o d e _ x o r :           s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 0 0 0 " ;               - -   0 x 0  
         c o n s t a n t   o p c o d e _ s e q :           s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 0 0 0 " ;               - -   0 x 0  
         c o n s t a n t   o p c o d e _ s n e :           s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 0 0 0 " ;               - -   0 x 0  
         c o n s t a n t   o p c o d e _ s l t :           s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 0 0 0 " ;               - -   0 x 0  
         c o n s t a n t   o p c o d e _ s g t :           s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 0 0 0 " ;               - -   0 x 0  
         c o n s t a n t   o p c o d e _ s l e :           s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 0 0 0 " ;               - -   0 x 0  
         c o n s t a n t   o p c o d e _ s g e :           s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 0 0 0 " ;               - -   0 x 0  
         c o n s t a n t   o p c o d e _ m o v i 2 s :     s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 0 0 0 " ;               - -   0 x 0  
         c o n s t a n t   o p c o d e _ m o v s 2 i :     s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 0 0 0 " ;               - -   0 x 0  
         c o n s t a n t   o p c o d e _ m o v f :         s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 0 0 0 " ;               - -   0 x 0  
         c o n s t a n t   o p c o d e _ m o v d :         s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 0 0 0 " ;               - -   0 x 0  
         c o n s t a n t   o p c o d e _ m o v f p 2 i :   s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 0 0 0 " ;               - -   0 x 0  
         c o n s t a n t   o p c o d e _ m o v i 2 f p :   s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 0 0 0 " ;               - -   0 x 0  
         c o n s t a n t   o p c o d e _ m o v i 2 t :     s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 0 0 0 " ;               - -   0 x 0  
         c o n s t a n t   o p c o d e _ m o v t 2 i :     s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 0 0 0 " ;               - -   0 x 0  
         c o n s t a n t   o p c o d e _ s l t u :         s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 0 0 0 " ;               - -   0 x 0  
         c o n s t a n t   o p c o d e _ s g t u :         s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 0 0 0 " ;               - -   0 x 0  
         c o n s t a n t   o p c o d e _ s l e u :         s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 0 0 0 " ;               - -   0 x 0  
         c o n s t a n t   o p c o d e _ s g e u :         s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 0 0 0 " ;               - -   0 x 0  
         c o n s t a n t   o p c o d e _ a d d f :         s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 1 0 0 " ;               - -   0 x 4  
         c o n s t a n t   o p c o d e _ s u b f :         s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 1 0 0 " ;               - -   0 x 4  
         c o n s t a n t   o p c o d e _ m u l t f :       s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 1 0 0 " ;               - -   0 x 4  
         c o n s t a n t   o p c o d e _ d i v f :         s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 1 0 0 " ;               - -   0 x 4  
         c o n s t a n t   o p c o d e _ a d d d :         s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 1 0 0 " ;               - -   0 x 4  
         c o n s t a n t   o p c o d e _ s u b d :         s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 1 0 0 " ;               - -   0 x 4  
         c o n s t a n t   o p c o d e _ m u l t d :       s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 1 0 0 " ;               - -   0 x 4  
         c o n s t a n t   o p c o d e _ d i v d :         s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 1 0 0 " ;               - -   0 x 4  
         c o n s t a n t   o p c o d e _ c v t f 2 d :     s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 1 0 0 " ;               - -   0 x 4  
         c o n s t a n t   o p c o d e _ c v t f 2 i :     s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 1 0 0 " ;               - -   0 x 4  
         c o n s t a n t   o p c o d e _ c v t d 2 f :     s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 1 0 0 " ;               - -   0 x 4  
         c o n s t a n t   o p c o d e _ c v t d 2 i :     s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 1 0 0 " ;               - -   0 x 4  
         c o n s t a n t   o p c o d e _ c v t i 2 f :     s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 1 0 0 " ;               - -   0 x 4  
         c o n s t a n t   o p c o d e _ c v t i 2 d :     s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 1 0 0 " ;               - -   0 x 4  
         c o n s t a n t   o p c o d e _ m u l t :         s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 1 0 0 " ;               - -   0 x 4  
         c o n s t a n t   o p c o d e _ d i v :           s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 1 0 0 " ;               - -   0 x 4  
         c o n s t a n t   o p c o d e _ e q f :           s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 1 0 0 " ;               - -   0 x 4  
         c o n s t a n t   o p c o d e _ n e f :           s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 1 0 0 " ;               - -   0 x 4  
         c o n s t a n t   o p c o d e _ l t f :           s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 1 0 0 " ;               - -   0 x 4  
         c o n s t a n t   o p c o d e _ g t f :           s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 1 0 0 " ;               - -   0 x 4  
         c o n s t a n t   o p c o d e _ l e f :           s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 1 0 0 " ;               - -   0 x 4  
         c o n s t a n t   o p c o d e _ g e f :           s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 1 0 0 " ;               - -   0 x 4  
         c o n s t a n t   o p c o d e _ m u l t u :       s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 1 0 0 " ;               - -   0 x 4  
         c o n s t a n t   o p c o d e _ d i v u :         s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 1 0 0 " ;               - -   0 x 4  
         c o n s t a n t   o p c o d e _ e q d :           s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 1 0 0 " ;               - -   0 x 4  
         c o n s t a n t   o p c o d e _ n e d :           s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 1 0 0 " ;               - -   0 x 4  
         c o n s t a n t   o p c o d e _ l t d :           s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 1 0 0 " ;               - -   0 x 4  
         c o n s t a n t   o p c o d e _ g t d :           s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 1 0 0 " ;               - -   0 x 4  
         c o n s t a n t   o p c o d e _ l e d :           s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 1 0 0 " ;               - -   0 x 4  
         c o n s t a n t   o p c o d e _ g e d :           s t d _ l o g i c _ v e c t o r ( 5   d o w n t o   0 )   : =   " 0 0 0 1 0 0 " ;               - -   0 x 4  
  
         - -   F U N C   F I E L D  
         c o n s t a n t   f u n c _ s l l :               s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 0 0 0 1 0 0 " ;   - -   0 x 0 4  
         c o n s t a n t   f u n c _ s r l :               s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 0 0 0 1 1 0 " ;   - -   0 x 0 6  
         c o n s t a n t   f u n c _ s r a :               s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 0 0 0 1 1 1 " ;   - -   0 x 0 7  
         c o n s t a n t   f u n c _ a d d :               s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 1 0 0 0 0 0 " ;   - -   0 x 2 0  
         c o n s t a n t   f u n c _ a d d u :             s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 1 0 0 0 0 1 " ;   - -   0 x 2 1  
         c o n s t a n t   f u n c _ s u b :               s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 1 0 0 0 1 0 " ;   - -   0 x 2 2  
         c o n s t a n t   f u n c _ s u b u :             s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 1 0 0 0 1 1 " ;   - -   0 x 2 3  
         c o n s t a n t   f u n c _ a n d :               s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 1 0 0 1 0 0 " ;   - -   0 x 2 4  
         c o n s t a n t   f u n c _ o r :                 s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 1 0 0 1 0 1 " ;   - -   0 x 2 5  
         c o n s t a n t   f u n c _ x o r :               s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 1 0 0 1 1 0 " ;   - -   0 x 2 6  
         c o n s t a n t   f u n c _ s e q :               s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 1 0 1 0 0 0 " ;   - -   0 x 2 8  
         c o n s t a n t   f u n c _ s n e :               s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 1 0 1 0 0 1 " ;   - -   0 x 2 9  
         c o n s t a n t   f u n c _ s l t :               s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 1 0 1 0 1 0 " ;   - -   0 x 2 a  
         c o n s t a n t   f u n c _ s g t :               s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 1 0 1 0 1 1 " ;   - -   0 x 2 b  
         c o n s t a n t   f u n c _ s l e :               s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 1 0 1 1 0 0 " ;   - -   0 x 2 c  
         c o n s t a n t   f u n c _ s g e :               s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 1 0 1 1 0 1 " ;   - -   0 x 2 d  
         c o n s t a n t   f u n c _ m o v i 2 s :         s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 1 1 0 0 0 0 " ;   - -   0 x 3 0  
         c o n s t a n t   f u n c _ m o v s 2 i :         s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 1 1 0 0 0 1 " ;   - -   0 x 3 1  
         c o n s t a n t   f u n c _ m o v f :             s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 1 1 0 0 1 0 " ;   - -   0 x 3 2  
         c o n s t a n t   f u n c _ m o v d :             s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 1 1 0 0 1 1 " ;   - -   0 x 3 3  
         c o n s t a n t   f u n c _ m o v f p 2 i :       s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 1 1 0 1 0 0 " ;   - -   0 x 3 4  
         c o n s t a n t   f u n c _ m o v i 2 f p :       s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 1 1 0 1 0 1 " ;   - -   0 x 3 5  
         c o n s t a n t   f u n c _ m o v i 2 t :         s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 1 1 0 1 1 0 " ;   - -   0 x 3 6  
         c o n s t a n t   f u n c _ m o v t 2 i :         s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 1 1 0 1 1 1 " ;   - -   0 x 3 7  
         c o n s t a n t   f u n c _ s l t u :             s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 1 1 1 0 1 0 " ;   - -   0 x 3 a  
         c o n s t a n t   f u n c _ s g t u :             s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 1 1 1 0 1 1 " ;   - -   0 x 3 b  
         c o n s t a n t   f u n c _ s l e u :             s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 1 1 1 1 0 0 " ;   - -   0 x 3 c  
         c o n s t a n t   f u n c _ s g e u :             s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 1 1 1 1 0 1 " ;   - -   0 x 3 d  
         c o n s t a n t   f u n c _ a d d f :             s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 0 0 0 0 0 0 " ;   - -   0 x 0 0  
         c o n s t a n t   f u n c _ s u b f :             s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 0 0 0 0 0 1 " ;   - -   0 x 0 1  
         c o n s t a n t   f u n c _ m u l t f :           s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 0 0 0 0 1 0 " ;   - -   0 x 0 2  
         c o n s t a n t   f u n c _ d i v f :             s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 0 0 0 0 1 1 " ;   - -   0 x 0 3  
         c o n s t a n t   f u n c _ a d d d :             s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 0 0 0 1 0 0 " ;   - -   0 x 0 4  
         c o n s t a n t   f u n c _ s u b d :             s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 0 0 0 1 0 1 " ;   - -   0 x 0 5  
         c o n s t a n t   f u n c _ m u l t d :           s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 0 0 0 1 1 0 " ;   - -   0 x 0 6  
         c o n s t a n t   f u n c _ d i v d :             s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 0 0 0 1 1 1 " ;   - -   0 x 0 7  
         c o n s t a n t   f u n c _ c v t f 2 d :         s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 0 0 1 0 0 0 " ;   - -   0 x 0 8  
         c o n s t a n t   f u n c _ c v t f 2 i :         s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 0 0 1 0 0 1 " ;   - -   0 x 0 9  
         c o n s t a n t   f u n c _ c v t d 2 f :         s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 0 0 1 0 1 0 " ;   - -   0 x 0 a  
         c o n s t a n t   f u n c _ c v t d 2 i :         s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 0 0 1 0 1 1 " ;   - -   0 x 0 b  
         c o n s t a n t   f u n c _ c v t i 2 f :         s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 0 0 1 1 0 0 " ;   - -   0 x 0 c  
         c o n s t a n t   f u n c _ c v t i 2 d :         s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 0 0 1 1 0 1 " ;   - -   0 x 0 d  
         c o n s t a n t   f u n c _ m u l t :             s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 0 0 1 1 1 0 " ;   - -   0 x 0 e  
         c o n s t a n t   f u n c _ d i v :               s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 0 0 1 1 1 1 " ;   - -   0 x 0 f  
         c o n s t a n t   f u n c _ e q f :               s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 0 1 0 0 0 0 " ;   - -   0 x 1 0  
         c o n s t a n t   f u n c _ n e f :               s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 0 1 0 0 0 1 " ;   - -   0 x 1 1  
         c o n s t a n t   f u n c _ l t f :               s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 0 1 0 0 1 0 " ;   - -   0 x 1 2  
         c o n s t a n t   f u n c _ g t f :               s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 0 1 0 0 1 1 " ;   - -   0 x 1 3  
         c o n s t a n t   f u n c _ l e f :               s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 0 1 0 1 0 0 " ;   - -   0 x 1 4  
         c o n s t a n t   f u n c _ g e f :               s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 0 1 0 1 0 1 " ;   - -   0 x 1 5  
         c o n s t a n t   f u n c _ m u l t u :           s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 0 1 0 1 1 0 " ;   - -   0 x 1 6  
         c o n s t a n t   f u n c _ d i v u :             s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 0 1 0 1 1 1 " ;   - -   0 x 1 7  
         c o n s t a n t   f u n c _ e q d :               s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 0 1 1 0 0 0 " ;   - -   0 x 1 8  
         c o n s t a n t   f u n c _ n e d :               s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 0 1 1 0 0 1 " ;   - -   0 x 1 9  
         c o n s t a n t   f u n c _ l t d :               s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 0 1 1 0 1 0 " ;   - -   0 x 1 a  
         c o n s t a n t   f u n c _ g t d :               s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 0 1 1 0 1 1 " ;   - -   0 x 1 b  
         c o n s t a n t   f u n c _ l e d :               s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 0 1 1 1 0 0 " ;   - -   0 x 1 c  
         c o n s t a n t   f u n c _ g e d :               s t d _ l o g i c _ v e c t o r ( 1 0   d o w n t o   0 )   : =   " 0 0 0 0 0 0 1 1 1 0 1 " ;   - -   0 x 1 d  
 e n d   i n s t r u c t i o n s _ p k g ;  
 